
module embedded_system (
	clk_clk,
	to_hex_readdata,
	reset_reset_n);	

	input		clk_clk;
	output	[31:0]	to_hex_readdata;
	input		reset_reset_n;
endmodule
