
module issp_test (
	source,
	probe);	

	output	[1:0]	source;
	input	[1:0]	probe;
endmodule
