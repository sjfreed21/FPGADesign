`ifdef sixforty
    parameter hArea = 800;
    parameter hFPorch = 16;
    parameter hBPorch = 48;
    parameter hSTime = 96;
    parameter vArea = 525;
    parameter vFPorch = 10;
    parameter vBPorch = 33;
    parameter vSTime = 2;
`endif