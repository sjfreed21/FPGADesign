parameter RESET = 4'b0000;
parameter START = 4'b0001;
parameter SENDA = 4'b0010;
parameter ACK_1 = 4'b0011;
parameter SEND1 = 4'b0100;
parameter ACK_2 = 4'b0101;
parameter SEND2 = 4'b0110;
parameter ACK_3 = 4'b0111;
parameter STOPC = 4'b1000;