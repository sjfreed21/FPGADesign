module pg(
    input  [9:0] hPixel,
    input  [8:0] vLine,
    input  [9:0] SW,
    output [7:0] RED,
    output [7:0] GRN,
    output [7:0] BLU
);